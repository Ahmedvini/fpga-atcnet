mirallll