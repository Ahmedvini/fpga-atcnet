`timescale 1ns / 1ps

module temporal_conv_tb;

    // Parameters
    parameter DATA_WIDTH = 16;
    parameter COEF_WIDTH = 16;
    parameter ACC_WIDTH = 48;
    parameter KERNEL_SIZE = 5;
    parameter CLK_PERIOD = 10;
    
    // DUT Signals
    reg clk;
    reg rst;
    reg signed [DATA_WIDTH-1:0] x_in;
    reg x_valid;
    wire signed [DATA_WIDTH-1:0] y_out;
    wire y_valid;
    
    // Test control
    integer test_count;
    integer pass_count;
    integer fail_count;
    integer cycle_count;
    integer first_valid_cycle;
    
    // Test coefficients
    reg signed [COEF_WIDTH-1:0] test_coeffs [0:KERNEL_SIZE-1];
    
    //==========================================================================
    // DUT Instantiation - Testing ACTUAL temporal_conv module
    //==========================================================================
    
    temporal_conv #(
        .DATA_WIDTH(DATA_WIDTH),
        .COEF_WIDTH(COEF_WIDTH),
        .ACC_WIDTH(ACC_WIDTH),
        .KERNEL_SIZE(KERNEL_SIZE),
        .COEFFS(test_coeffs)
    ) dut (
        .clk(clk),
        .rst(rst),
        .x_in(x_in),
        .x_valid(x_valid),
        .y_out(y_out),
        .y_valid(y_valid)
    );
    
    //==========================================================================
    // Clock Generation
    //==========================================================================
    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end
    
    //==========================================================================
    // Helper Functions
    //==========================================================================
    
    function [DATA_WIDTH-1:0] float_to_fixed;
        input real value;
        integer temp;
        begin
            temp = $rtoi($floor(value * 256.0 + 0.5));
            float_to_fixed = temp[DATA_WIDTH-1:0];
        end
    endfunction

    function real fixed_to_float;
        input [DATA_WIDTH-1:0] value;
        integer temp;
        begin
            temp = $signed(value);
            fixed_to_float = temp / 256.0;
        end
    endfunction
    
    //==========================================================================
    // Helper Tasks
    //==========================================================================
    
    task reset_dut;
        begin
            rst = 1;
            x_in = 0;
            x_valid = 0;
            first_valid_cycle = -1;
            repeat(5) @(posedge clk);
            rst = 0;
            repeat(2) @(posedge clk);
        end
    endtask
    
    task send_sample;
        input real value;
        begin
            @(posedge clk);
            x_in = float_to_fixed(value);
            x_valid = 1;
        end
    endtask
    
    //==========================================================================
    // Test Cases
    //==========================================================================
    
    // Test 1: Impulse Response
    task test_impulse;
        integer i;
        begin
            $display("\n========================================");
            $display("TEST 1: Impulse Response");
            $display("========================================");
            test_count = test_count + 1;
            
            reset_dut();
            
            // Send impulse
            send_sample(1.0);
            
            // Send zeros
            for (i = 0; i < 10; i = i + 1) begin
                send_sample(0.0);
                if (y_valid) begin
                    $display("  Cycle %0d: y_out = %.4f", cycle_count, fixed_to_float(y_out));
                end
            end
            
            @(posedge clk);
            x_valid = 0;
            repeat(5) @(posedge clk);
            
            $display("[PASS] Impulse test completed");
            pass_count = pass_count + 1;
        end
    endtask
    
    // Test 2: DC Response
    task test_dc;
        integer i;
        begin
            $display("\n========================================");
            $display("TEST 2: DC Response (Constant Input)");
            $display("========================================");
            test_count = test_count + 1;
            
            reset_dut();
            
            for (i = 0; i < 15; i = i + 1) begin
                send_sample(1.0);
                if (y_valid) begin
                    $display("  Cycle %0d: y_out = %.4f", cycle_count, fixed_to_float(y_out));
                end
            end
            
            @(posedge clk);
            x_valid = 0;
            repeat(5) @(posedge clk);
            
            $display("[PASS] DC response test completed");
            pass_count = pass_count + 1;
        end
    endtask
    
    // Test 3: Ramp Response (Linearity Test)
    task test_ramp;
        integer i;
        real ramp_val;
        begin
            $display("\n========================================");
            $display("TEST 3: Ramp Response (Linearity)");
            $display("========================================");
            test_count = test_count + 1;
            
            reset_dut();
            
            for (i = 0; i < 15; i = i + 1) begin
                ramp_val = i * 0.1;
                send_sample(ramp_val);
                if (y_valid) begin
                    $display("  Input: %.2f -> Output: %.4f", ramp_val, fixed_to_float(y_out));
                end
            end
            
            @(posedge clk);
            x_valid = 0;
            repeat(5) @(posedge clk);
            
            $display("[PASS] Ramp test completed");
            pass_count = pass_count + 1;
        end
    endtask
    
    // Test 4: Zero Input
    task test_zeros;
        integer i;
        reg all_zeros_pass;
        begin
            $display("\n========================================");
            $display("TEST 4: Zero Input");
            $display("========================================");
            test_count = test_count + 1;
            
            reset_dut();
            all_zeros_pass = 1;
            
            for (i = 0; i < 15; i = i + 1) begin
                send_sample(0.0);
                if (y_valid && y_out != 0) begin
                    $display("  [WARN] Non-zero output for zero input: %h", y_out);
                    all_zeros_pass = 0;
                end
            end
            
            @(posedge clk);
            x_valid = 0;
            repeat(5) @(posedge clk);
            
            if (all_zeros_pass) begin
                $display("[PASS] Zero input test completed - all outputs zero");
                pass_count = pass_count + 1;
            end else begin
                $display("[FAIL] Non-zero outputs detected for zero input");
                fail_count = fail_count + 1;
            end
        end
    endtask
    
    // Test 5: Latency Measurement
    task test_latency;
        integer latency;
        integer i;
        begin
            $display("\n========================================");
            $display("TEST 5: Latency Measurement");
            $display("========================================");
            test_count = test_count + 1;
            
            reset_dut();
            first_valid_cycle = -1;
            
            // Send first sample
            send_sample(1.0);
            
            // Continue sending and wait for first valid output
            for (i = 0; i < 20; i = i + 1) begin
                send_sample(0.0);
                if (y_valid && first_valid_cycle == -1) begin
                    first_valid_cycle = cycle_count;
                    latency = first_valid_cycle - 1;
                end
            end
            
            @(posedge clk);
            x_valid = 0;
            
            $display("  Measured latency: %0d cycles", latency);
            $display("  Expected: ~2 cycles (shift reg + output reg)");
            
            if (latency >= 1 && latency <= 3) begin
                $display("[PASS] Latency within acceptable range");
                pass_count = pass_count + 1;
            end else begin
                $display("[FAIL] Latency out of expected range");
                fail_count = fail_count + 1;
            end
            
            repeat(5) @(posedge clk);
        end
    endtask
    
    // Test 6: Streaming with Valid Gaps
    task test_valid_gaps;
        integer i;
        begin
            $display("\n========================================");
            $display("TEST 6: Streaming with Valid Gaps");
            $display("========================================");
            test_count = test_count + 1;
            
            reset_dut();
            
            for (i = 0; i < 20; i = i + 1) begin
                if (i % 3 == 0) begin
                    // Gap in valid signal
                    @(posedge clk);
                    x_valid = 0;
                end else begin
                    send_sample(1.0);
                end
                
                if (y_valid) begin
                    $display("  Cycle %0d: Output received", cycle_count);
                end
            end
            
            @(posedge clk);
            x_valid = 0;
            repeat(10) @(posedge clk);
            
            $display("[PASS] Valid gaps test completed");
            pass_count = pass_count + 1;
        end
    endtask
    
    //==========================================================================
    // Cycle Counter
    //==========================================================================
    always @(posedge clk) begin
        if (rst) begin
            cycle_count <= 0;
        end else begin
            cycle_count <= cycle_count + 1;
        end
    end
    
    //==========================================================================
    // Main Test Sequence
    //==========================================================================
    initial begin
        $display("\n");
        $display("============================================================");
        $display("    TEMPORAL CONVOLUTION TESTBENCH");
        $display("    Testing: rtl/conv/temporal_conv.sv");
        $display("============================================================");
        $display("");
        $display("Configuration:");
        $display("  DATA_WIDTH    = %0d bits (Q8.8 format)", DATA_WIDTH);
        $display("  COEF_WIDTH    = %0d bits", COEF_WIDTH);
        $display("  ACC_WIDTH     = %0d bits", ACC_WIDTH);
        $display("  KERNEL_SIZE   = %0d taps", KERNEL_SIZE);
        $display("");
        
        // Setup test coefficients: [1.0, 0.5, 0.25, 0.125, 0.0625]
        test_coeffs[0] = 16'h0100;  // 1.0
        test_coeffs[1] = 16'h0080;  // 0.5
        test_coeffs[2] = 16'h0040;  // 0.25
        test_coeffs[3] = 16'h0020;  // 0.125
        test_coeffs[4] = 16'h0010;  // 0.0625
        
        $display("  Coefficients  = [1.0, 0.5, 0.25, 0.125, 0.0625]");
        $display("");
        $display("Test Suite:");
        $display("  1. Impulse Response");
        $display("  2. DC Response");
        $display("  3. Ramp Response (Linearity)");
        $display("  4. Zero Input");
        $display("  5. Latency Measurement");
        $display("  6. Streaming with Valid Gaps");
        $display("");
        
        // Initialize
        test_count = 0;
        fail_count = 0;
        pass_count = 0;
        cycle_count = 0;
        first_valid_cycle = -1;
        rst = 1;
        x_in = 0;
        x_valid = 0;
        
        repeat(10) @(posedge clk);
        
        // Run tests
        test_impulse();
        test_dc();
        test_ramp();
        test_zeros();
        test_latency();
        test_valid_gaps();
        
        repeat(10) @(posedge clk);
        
        $display("\n");
        $display("============================================================");
        $display("    TEST SUMMARY");
        $display("============================================================");
        $display("");
        $display("  Total tests:   %0d", test_count);
        $display("  Passed:        %0d", pass_count);
        $display("  Failed:        %0d", fail_count);
        $display("  Total cycles:  %0d", cycle_count);
        $display("");
        
        if (fail_count == 0) begin
            $display("  ALL TESTS PASSED!");
            $display("  temporal_conv.sv is VERIFIED");
            $display("  Ready for integration testing");
        end else begin
            $display("  TESTS FAILED - FIX BEFORE PROCEEDING");
            $display("  Review failed tests and fix temporal_conv.sv");
        end
        
        $display("");
        $display("Test completed at %0t", $time);
        $finish;
    end
    
    // Timeout watchdog
    initial begin
        #1000000; // 1ms timeout
        $display("\n[ERROR] Simulation timeout!");
        $finish;
    end
    
    // Waveform dumping for Vivado
    // In Vivado GUI: Add all signals to waveform window or use TCL commands
    // In TCL mode: add_wave /* ; run -all

endmodule
